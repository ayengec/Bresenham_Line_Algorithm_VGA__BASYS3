package testbench_pkg;
   // `include "vga_interface.sv"
    `include "const_pkg.svh"
    `include "sequence_item.svh"
    `include "generator.svh"
    `include "driver.svh"
    `include "monitor.svh"
    `include "scoreboard.svh"
    `include "environment.svh"
    `include "test.svh"
endpackage